module not_5(out,in);

input [4:0]in;
output [4:0]out;
not (out[0],in[0]);
not (out[1],in[1]);
not (out[2],in[2]);
not (out[3],in[3]);
not (out[4],in[4]);
endmodule